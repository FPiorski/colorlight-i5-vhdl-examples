LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY character_ram IS
    GENERIC
    (
        g_depth_log2 : positive;
        g_char_w     : positive;
        g_char_h     : positive
    );
    PORT
    (
        i_clk        : IN    std_logic;

        i_wr_addr    : IN    std_logic_vector(g_depth_log2-1 downto 0);
        i_wr_data    : IN    std_logic_vector(    g_char_w-1 downto 0);
        i_wr_ena     : IN    std_logic;

        i_rd_addr    : IN    std_logic_vector(g_depth_log2-1 downto 0);
        o_rd_data    :   OUT std_logic_vector(    g_char_w-1 downto 0)
    );
END character_ram;

ARCHITECTURE RTL OF character_ram IS

    CONSTANT C_depth    : integer := 2**g_depth_log2;

    TYPE     T_char_arr IS ARRAY (0 TO C_depth-1) OF std_logic_vector(g_char_h-1 downto 0);

    FUNCTION f_init_char_arr RETURN T_char_arr is
        VARIABLE v_return    : T_char_arr := (OTHERS => (OTHERS => '0'));
    BEGIN
        IF (g_char_w = 8 AND g_char_h = 8) THEN
            REPORT "character_ram: 8x8 characters, initializing stored font";
            FOR code IN 0 TO 2**g_depth_log2-1 LOOP
                CASE code IS
                    WHEN 0 =>
                        v_return(code*g_char_h + 0) := "11110000";
                        v_return(code*g_char_h + 1) := "10010000";
                        v_return(code*g_char_h + 2) := "10010000";
                        v_return(code*g_char_h + 3) := "10010000";
                        v_return(code*g_char_h + 4) := "11110000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 1 =>
                        v_return(code*g_char_h + 0) := "01100000";
                        v_return(code*g_char_h + 1) := "10100000";
                        v_return(code*g_char_h + 2) := "00100000";
                        v_return(code*g_char_h + 3) := "00100000";
                        v_return(code*g_char_h + 4) := "11110000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 2 =>
                        v_return(code*g_char_h + 0) := "01100000";
                        v_return(code*g_char_h + 1) := "10010000";
                        v_return(code*g_char_h + 2) := "01100000";
                        v_return(code*g_char_h + 3) := "10000000";
                        v_return(code*g_char_h + 4) := "11110000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 3 =>
                        v_return(code*g_char_h + 0) := "11110000";
                        v_return(code*g_char_h + 1) := "00010000";
                        v_return(code*g_char_h + 2) := "11110000";
                        v_return(code*g_char_h + 3) := "00010000";
                        v_return(code*g_char_h + 4) := "11110000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 4 =>
                        v_return(code*g_char_h + 0) := "10000000";
                        v_return(code*g_char_h + 1) := "10000000";
                        v_return(code*g_char_h + 2) := "11110000";
                        v_return(code*g_char_h + 3) := "00100000";
                        v_return(code*g_char_h + 4) := "00100000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 5 =>
                        v_return(code*g_char_h + 0) := "11110000";
                        v_return(code*g_char_h + 1) := "10000000";
                        v_return(code*g_char_h + 2) := "11100000";
                        v_return(code*g_char_h + 3) := "00010000";
                        v_return(code*g_char_h + 4) := "11100000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 6 =>
                        v_return(code*g_char_h + 0) := "01110000";
                        v_return(code*g_char_h + 1) := "10000000";
                        v_return(code*g_char_h + 2) := "11100000";
                        v_return(code*g_char_h + 3) := "10010000";
                        v_return(code*g_char_h + 4) := "11100000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 7 =>
                        v_return(code*g_char_h + 0) := "11110000";
                        v_return(code*g_char_h + 1) := "00010000";
                        v_return(code*g_char_h + 2) := "00100000";
                        v_return(code*g_char_h + 3) := "01000000";
                        v_return(code*g_char_h + 4) := "10000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 8 =>
                        v_return(code*g_char_h + 0) := "01100000";
                        v_return(code*g_char_h + 1) := "10010000";
                        v_return(code*g_char_h + 2) := "01100000";
                        v_return(code*g_char_h + 3) := "10010000";
                        v_return(code*g_char_h + 4) := "01100000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 9 =>
                        v_return(code*g_char_h + 0) := "01100000";
                        v_return(code*g_char_h + 1) := "10010000";
                        v_return(code*g_char_h + 2) := "01110000";
                        v_return(code*g_char_h + 3) := "00010000";
                        v_return(code*g_char_h + 4) := "11100000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 10 =>
                        v_return(code*g_char_h + 0) := "01100000";
                        v_return(code*g_char_h + 1) := "10010000";
                        v_return(code*g_char_h + 2) := "11110000";
                        v_return(code*g_char_h + 3) := "10010000";
                        v_return(code*g_char_h + 4) := "10010000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 11 =>
                        v_return(code*g_char_h + 0) := "11100000";
                        v_return(code*g_char_h + 1) := "10010000";
                        v_return(code*g_char_h + 2) := "11100000";
                        v_return(code*g_char_h + 3) := "10010000";
                        v_return(code*g_char_h + 4) := "11100000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 12 =>
                        v_return(code*g_char_h + 0) := "01110000";
                        v_return(code*g_char_h + 1) := "10000000";
                        v_return(code*g_char_h + 2) := "10000000";
                        v_return(code*g_char_h + 3) := "10000000";
                        v_return(code*g_char_h + 4) := "01110000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 13 =>
                        v_return(code*g_char_h + 0) := "11100000";
                        v_return(code*g_char_h + 1) := "10010000";
                        v_return(code*g_char_h + 2) := "10010000";
                        v_return(code*g_char_h + 3) := "10010000";
                        v_return(code*g_char_h + 4) := "11100000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 14 =>
                        v_return(code*g_char_h + 0) := "11110000";
                        v_return(code*g_char_h + 1) := "10000000";
                        v_return(code*g_char_h + 2) := "11110000";
                        v_return(code*g_char_h + 3) := "10000000";
                        v_return(code*g_char_h + 4) := "11110000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 15 =>
                        v_return(code*g_char_h + 0) := "11110000";
                        v_return(code*g_char_h + 1) := "10000000";
                        v_return(code*g_char_h + 2) := "11100000";
                        v_return(code*g_char_h + 3) := "10000000";
                        v_return(code*g_char_h + 4) := "10000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 16 =>
                        v_return(code*g_char_h + 0) := "01101111";
                        v_return(code*g_char_h + 1) := "10101001";
                        v_return(code*g_char_h + 2) := "00101001";
                        v_return(code*g_char_h + 3) := "00101001";
                        v_return(code*g_char_h + 4) := "11111111";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 17 =>
                        v_return(code*g_char_h + 0) := "01100110";
                        v_return(code*g_char_h + 1) := "10101010";
                        v_return(code*g_char_h + 2) := "00100010";
                        v_return(code*g_char_h + 3) := "00100010";
                        v_return(code*g_char_h + 4) := "11111111";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 18 =>
                        v_return(code*g_char_h + 0) := "01100110";
                        v_return(code*g_char_h + 1) := "10101001";
                        v_return(code*g_char_h + 2) := "00100110";
                        v_return(code*g_char_h + 3) := "00101000";
                        v_return(code*g_char_h + 4) := "11111111";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 19 =>
                        v_return(code*g_char_h + 0) := "01101111";
                        v_return(code*g_char_h + 1) := "10100001";
                        v_return(code*g_char_h + 2) := "00101111";
                        v_return(code*g_char_h + 3) := "00100001";
                        v_return(code*g_char_h + 4) := "11111111";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 20 =>
                        v_return(code*g_char_h + 0) := "01101000";
                        v_return(code*g_char_h + 1) := "10101000";
                        v_return(code*g_char_h + 2) := "00101111";
                        v_return(code*g_char_h + 3) := "00100010";
                        v_return(code*g_char_h + 4) := "11110010";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 21 =>
                        v_return(code*g_char_h + 0) := "01101111";
                        v_return(code*g_char_h + 1) := "10101000";
                        v_return(code*g_char_h + 2) := "00101110";
                        v_return(code*g_char_h + 3) := "00100001";
                        v_return(code*g_char_h + 4) := "11111110";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 22 =>
                        v_return(code*g_char_h + 0) := "01100111";
                        v_return(code*g_char_h + 1) := "10101000";
                        v_return(code*g_char_h + 2) := "00101110";
                        v_return(code*g_char_h + 3) := "00101001";
                        v_return(code*g_char_h + 4) := "11111110";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 23 =>
                        v_return(code*g_char_h + 0) := "01101111";
                        v_return(code*g_char_h + 1) := "10100001";
                        v_return(code*g_char_h + 2) := "00100010";
                        v_return(code*g_char_h + 3) := "00100100";
                        v_return(code*g_char_h + 4) := "11111000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 24 =>
                        v_return(code*g_char_h + 0) := "01100110";
                        v_return(code*g_char_h + 1) := "10101001";
                        v_return(code*g_char_h + 2) := "00100110";
                        v_return(code*g_char_h + 3) := "00101001";
                        v_return(code*g_char_h + 4) := "11110110";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 25 =>
                        v_return(code*g_char_h + 0) := "01100110";
                        v_return(code*g_char_h + 1) := "10101001";
                        v_return(code*g_char_h + 2) := "00100111";
                        v_return(code*g_char_h + 3) := "00100001";
                        v_return(code*g_char_h + 4) := "11111110";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 26 =>
                        v_return(code*g_char_h + 0) := "01100110";
                        v_return(code*g_char_h + 1) := "10101001";
                        v_return(code*g_char_h + 2) := "00101111";
                        v_return(code*g_char_h + 3) := "00101001";
                        v_return(code*g_char_h + 4) := "11111001";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 27 =>
                        v_return(code*g_char_h + 0) := "01101110";
                        v_return(code*g_char_h + 1) := "10101001";
                        v_return(code*g_char_h + 2) := "00101110";
                        v_return(code*g_char_h + 3) := "00101001";
                        v_return(code*g_char_h + 4) := "11111110";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 28 =>
                        v_return(code*g_char_h + 0) := "01100111";
                        v_return(code*g_char_h + 1) := "10101000";
                        v_return(code*g_char_h + 2) := "00101000";
                        v_return(code*g_char_h + 3) := "00101000";
                        v_return(code*g_char_h + 4) := "11110111";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 29 =>
                        v_return(code*g_char_h + 0) := "01101110";
                        v_return(code*g_char_h + 1) := "10101001";
                        v_return(code*g_char_h + 2) := "00101001";
                        v_return(code*g_char_h + 3) := "00101001";
                        v_return(code*g_char_h + 4) := "11111110";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 30 =>
                        v_return(code*g_char_h + 0) := "01101111";
                        v_return(code*g_char_h + 1) := "10101000";
                        v_return(code*g_char_h + 2) := "00101111";
                        v_return(code*g_char_h + 3) := "00101000";
                        v_return(code*g_char_h + 4) := "11111111";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 31 =>
                        v_return(code*g_char_h + 0) := "01101111";
                        v_return(code*g_char_h + 1) := "10101000";
                        v_return(code*g_char_h + 2) := "00101110";
                        v_return(code*g_char_h + 3) := "00101000";
                        v_return(code*g_char_h + 4) := "11111000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 32 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 33 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00011000";
                        v_return(code*g_char_h + 2) := "00011000";
                        v_return(code*g_char_h + 3) := "00011000";
                        v_return(code*g_char_h + 4) := "00011000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00011000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 34 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "01100110";
                        v_return(code*g_char_h + 2) := "01100110";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 35 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00100100";
                        v_return(code*g_char_h + 2) := "01111110";
                        v_return(code*g_char_h + 3) := "00100100";
                        v_return(code*g_char_h + 4) := "00100100";
                        v_return(code*g_char_h + 5) := "01111110";
                        v_return(code*g_char_h + 6) := "00100100";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 36 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00001000";
                        v_return(code*g_char_h + 2) := "00111110";
                        v_return(code*g_char_h + 3) := "01001000";
                        v_return(code*g_char_h + 4) := "00111100";
                        v_return(code*g_char_h + 5) := "00001010";
                        v_return(code*g_char_h + 6) := "01111100";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 37 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 38 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 39 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 40 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 41 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 42 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"14";
                        v_return(code*g_char_h + 2) := X"08";
                        v_return(code*g_char_h + 3) := X"14";
                        v_return(code*g_char_h + 4) := X"00";
                        v_return(code*g_char_h + 5) := X"00";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 43 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"10";
                        v_return(code*g_char_h + 3) := X"38";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"00";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 44 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"00";
                        v_return(code*g_char_h + 3) := X"00";
                        v_return(code*g_char_h + 4) := X"00";
                        v_return(code*g_char_h + 5) := X"10";
                        v_return(code*g_char_h + 6) := X"10";
                        v_return(code*g_char_h + 7) := X"20";
                    WHEN 45 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"00";
                        v_return(code*g_char_h + 3) := X"3C";
                        v_return(code*g_char_h + 4) := X"00";
                        v_return(code*g_char_h + 5) := X"00";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 46 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"00";
                        v_return(code*g_char_h + 3) := X"00";
                        v_return(code*g_char_h + 4) := X"00";
                        v_return(code*g_char_h + 5) := X"08";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 47 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"02";
                        v_return(code*g_char_h + 2) := X"04";
                        v_return(code*g_char_h + 3) := X"08";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"20";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 48 =>
                        v_return(code*g_char_h + 0) := X"18";
                        v_return(code*g_char_h + 1) := X"24";
                        v_return(code*g_char_h + 2) := X"24";
                        v_return(code*g_char_h + 3) := X"24";
                        v_return(code*g_char_h + 4) := X"24";
                        v_return(code*g_char_h + 5) := X"18";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 49 =>
                        v_return(code*g_char_h + 0) := X"18";
                        v_return(code*g_char_h + 1) := X"28";
                        v_return(code*g_char_h + 2) := X"08";
                        v_return(code*g_char_h + 3) := X"08";
                        v_return(code*g_char_h + 4) := X"08";
                        v_return(code*g_char_h + 5) := X"3C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 50 =>
                        v_return(code*g_char_h + 0) := X"38";
                        v_return(code*g_char_h + 1) := X"44";
                        v_return(code*g_char_h + 2) := X"08";
                        v_return(code*g_char_h + 3) := X"10";
                        v_return(code*g_char_h + 4) := X"20";
                        v_return(code*g_char_h + 5) := X"7C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 51 =>
                        v_return(code*g_char_h + 0) := X"38";
                        v_return(code*g_char_h + 1) := X"44";
                        v_return(code*g_char_h + 2) := X"04";
                        v_return(code*g_char_h + 3) := X"18";
                        v_return(code*g_char_h + 4) := X"44";
                        v_return(code*g_char_h + 5) := X"38";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 52 =>
                        v_return(code*g_char_h + 0) := X"20";
                        v_return(code*g_char_h + 1) := X"20";
                        v_return(code*g_char_h + 2) := X"24";
                        v_return(code*g_char_h + 3) := X"3E";
                        v_return(code*g_char_h + 4) := X"04";
                        v_return(code*g_char_h + 5) := X"04";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 53 =>
                        v_return(code*g_char_h + 0) := X"3E";
                        v_return(code*g_char_h + 1) := X"20";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"02";
                        v_return(code*g_char_h + 4) := X"02";
                        v_return(code*g_char_h + 5) := X"3C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 54 =>
                        v_return(code*g_char_h + 0) := X"1C";
                        v_return(code*g_char_h + 1) := X"20";
                        v_return(code*g_char_h + 2) := X"38";
                        v_return(code*g_char_h + 3) := X"24";
                        v_return(code*g_char_h + 4) := X"24";
                        v_return(code*g_char_h + 5) := X"18";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 55 =>
                        v_return(code*g_char_h + 0) := X"3C";
                        v_return(code*g_char_h + 1) := X"44";
                        v_return(code*g_char_h + 2) := X"08";
                        v_return(code*g_char_h + 3) := X"10";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"10";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 56 =>
                        v_return(code*g_char_h + 0) := X"18";
                        v_return(code*g_char_h + 1) := X"24";
                        v_return(code*g_char_h + 2) := X"18";
                        v_return(code*g_char_h + 3) := X"24";
                        v_return(code*g_char_h + 4) := X"24";
                        v_return(code*g_char_h + 5) := X"18";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 57 =>
                        v_return(code*g_char_h + 0) := X"18";
                        v_return(code*g_char_h + 1) := X"24";
                        v_return(code*g_char_h + 2) := X"1C";
                        v_return(code*g_char_h + 3) := X"04";
                        v_return(code*g_char_h + 4) := X"04";
                        v_return(code*g_char_h + 5) := X"18";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 58 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"08";
                        v_return(code*g_char_h + 3) := X"00";
                        v_return(code*g_char_h + 4) := X"00";
                        v_return(code*g_char_h + 5) := X"08";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 59 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 60 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 61 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"00";
                        v_return(code*g_char_h + 4) := X"3C";
                        v_return(code*g_char_h + 5) := X"00";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 62 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 63 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 64 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 65 =>
                        v_return(code*g_char_h + 0) := X"18";
                        v_return(code*g_char_h + 1) := X"24";
                        v_return(code*g_char_h + 2) := X"24";
                        v_return(code*g_char_h + 3) := X"7E";
                        v_return(code*g_char_h + 4) := X"42";
                        v_return(code*g_char_h + 5) := X"42";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 66 =>
                        v_return(code*g_char_h + 0) := X"7C";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"7C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 67 =>
                        v_return(code*g_char_h + 0) := X"3C";
                        v_return(code*g_char_h + 1) := X"42";
                        v_return(code*g_char_h + 2) := X"40";
                        v_return(code*g_char_h + 3) := X"40";
                        v_return(code*g_char_h + 4) := X"42";
                        v_return(code*g_char_h + 5) := X"3C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 68 =>
                        v_return(code*g_char_h + 0) := X"7C";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"22";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"7C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 69 =>
                        v_return(code*g_char_h + 0) := X"7E";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"38";
                        v_return(code*g_char_h + 3) := X"20";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"7E";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 70 =>
                        v_return(code*g_char_h + 0) := X"7E";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"38";
                        v_return(code*g_char_h + 3) := X"20";
                        v_return(code*g_char_h + 4) := X"20";
                        v_return(code*g_char_h + 5) := X"70";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 71 =>
                        v_return(code*g_char_h + 0) := X"1C";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"20";
                        v_return(code*g_char_h + 3) := X"26";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"1C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 72 =>
                        v_return(code*g_char_h + 0) := X"44";
                        v_return(code*g_char_h + 1) := X"44";
                        v_return(code*g_char_h + 2) := X"7C";
                        v_return(code*g_char_h + 3) := X"44";
                        v_return(code*g_char_h + 4) := X"44";
                        v_return(code*g_char_h + 5) := X"44";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 73 =>
                        v_return(code*g_char_h + 0) := X"38";
                        v_return(code*g_char_h + 1) := X"10";
                        v_return(code*g_char_h + 2) := X"10";
                        v_return(code*g_char_h + 3) := X"10";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"38";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 74 =>
                        v_return(code*g_char_h + 0) := X"70";
                        v_return(code*g_char_h + 1) := X"10";
                        v_return(code*g_char_h + 2) := X"10";
                        v_return(code*g_char_h + 3) := X"90";
                        v_return(code*g_char_h + 4) := X"90";
                        v_return(code*g_char_h + 5) := X"70";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 75 =>
                        v_return(code*g_char_h + 0) := X"64";
                        v_return(code*g_char_h + 1) := X"28";
                        v_return(code*g_char_h + 2) := X"30";
                        v_return(code*g_char_h + 3) := X"28";
                        v_return(code*g_char_h + 4) := X"24";
                        v_return(code*g_char_h + 5) := X"64";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 76 =>
                        v_return(code*g_char_h + 0) := X"38";
                        v_return(code*g_char_h + 1) := X"10";
                        v_return(code*g_char_h + 2) := X"10";
                        v_return(code*g_char_h + 3) := X"10";
                        v_return(code*g_char_h + 4) := X"12";
                        v_return(code*g_char_h + 5) := X"1E";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 77 =>
                        v_return(code*g_char_h + 0) := X"22";
                        v_return(code*g_char_h + 1) := X"36";
                        v_return(code*g_char_h + 2) := X"2A";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"22";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 78 =>
                        v_return(code*g_char_h + 0) := X"22";
                        v_return(code*g_char_h + 1) := X"32";
                        v_return(code*g_char_h + 2) := X"2A";
                        v_return(code*g_char_h + 3) := X"26";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"22";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 79 =>
                        v_return(code*g_char_h + 0) := X"38";
                        v_return(code*g_char_h + 1) := X"44";
                        v_return(code*g_char_h + 2) := X"44";
                        v_return(code*g_char_h + 3) := X"44";
                        v_return(code*g_char_h + 4) := X"44";
                        v_return(code*g_char_h + 5) := X"38";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 80 =>
                        v_return(code*g_char_h + 0) := X"7C";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"20";
                        v_return(code*g_char_h + 4) := X"20";
                        v_return(code*g_char_h + 5) := X"70";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 81 =>
                        v_return(code*g_char_h + 0) := X"38";
                        v_return(code*g_char_h + 1) := X"44";
                        v_return(code*g_char_h + 2) := X"44";
                        v_return(code*g_char_h + 3) := X"44";
                        v_return(code*g_char_h + 4) := X"4C";
                        v_return(code*g_char_h + 5) := X"38";
                        v_return(code*g_char_h + 6) := X"08";
                        v_return(code*g_char_h + 7) := X"04";
                    WHEN 82 =>
                        v_return(code*g_char_h + 0) := X"7C";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"62";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 83 =>
                        v_return(code*g_char_h + 0) := X"18";
                        v_return(code*g_char_h + 1) := X"24";
                        v_return(code*g_char_h + 2) := X"10";
                        v_return(code*g_char_h + 3) := X"08";
                        v_return(code*g_char_h + 4) := X"24";
                        v_return(code*g_char_h + 5) := X"18";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 84 =>
                        v_return(code*g_char_h + 0) := X"7F";
                        v_return(code*g_char_h + 1) := X"49";
                        v_return(code*g_char_h + 2) := X"08";
                        v_return(code*g_char_h + 3) := X"08";
                        v_return(code*g_char_h + 4) := X"08";
                        v_return(code*g_char_h + 5) := X"1C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 85 =>
                        v_return(code*g_char_h + 0) := X"22";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"22";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"1C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 86 =>
                        v_return(code*g_char_h + 0) := X"22";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"22";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"14";
                        v_return(code*g_char_h + 5) := X"08";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 87 =>
                        v_return(code*g_char_h + 0) := X"22";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"22";
                        v_return(code*g_char_h + 3) := X"2A";
                        v_return(code*g_char_h + 4) := X"36";
                        v_return(code*g_char_h + 5) := X"22";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 88 =>
                        v_return(code*g_char_h + 0) := X"22";
                        v_return(code*g_char_h + 1) := X"14";
                        v_return(code*g_char_h + 2) := X"08";
                        v_return(code*g_char_h + 3) := X"14";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"22";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 89 =>
                        v_return(code*g_char_h + 0) := X"22";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"14";
                        v_return(code*g_char_h + 3) := X"08";
                        v_return(code*g_char_h + 4) := X"08";
                        v_return(code*g_char_h + 5) := X"1C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 90 =>
                        v_return(code*g_char_h + 0) := X"3E";
                        v_return(code*g_char_h + 1) := X"22";
                        v_return(code*g_char_h + 2) := X"04";
                        v_return(code*g_char_h + 3) := X"08";
                        v_return(code*g_char_h + 4) := X"12";
                        v_return(code*g_char_h + 5) := X"3E";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 91 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 92 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 93 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 94 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 95 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"00";
                        v_return(code*g_char_h + 3) := X"00";
                        v_return(code*g_char_h + 4) := X"00";
                        v_return(code*g_char_h + 5) := X"7E";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 96 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 97 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"38";
                        v_return(code*g_char_h + 3) := X"44";
                        v_return(code*g_char_h + 4) := X"44";
                        v_return(code*g_char_h + 5) := X"3E";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 98 =>
                        v_return(code*g_char_h + 0) := X"20";
                        v_return(code*g_char_h + 1) := X"20";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"3C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 99 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"1C";
                        v_return(code*g_char_h + 3) := X"20";
                        v_return(code*g_char_h + 4) := X"20";
                        v_return(code*g_char_h + 5) := X"1C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 100 =>
                        v_return(code*g_char_h + 0) := X"02";
                        v_return(code*g_char_h + 1) := X"02";
                        v_return(code*g_char_h + 2) := X"1E";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"1E";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 101 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"1C";
                        v_return(code*g_char_h + 2) := X"22";
                        v_return(code*g_char_h + 3) := X"3E";
                        v_return(code*g_char_h + 4) := X"20";
                        v_return(code*g_char_h + 5) := X"1C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 102 =>
                        v_return(code*g_char_h + 0) := X"18";
                        v_return(code*g_char_h + 1) := X"24";
                        v_return(code*g_char_h + 2) := X"20";
                        v_return(code*g_char_h + 3) := X"70";
                        v_return(code*g_char_h + 4) := X"20";
                        v_return(code*g_char_h + 5) := X"20";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 103 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"1C";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"1E";
                        v_return(code*g_char_h + 6) := X"02";
                        v_return(code*g_char_h + 7) := X"1C";
                    WHEN 104 =>
                        v_return(code*g_char_h + 0) := X"20";
                        v_return(code*g_char_h + 1) := X"20";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"22";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 105 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"10";
                        v_return(code*g_char_h + 2) := X"00";
                        v_return(code*g_char_h + 3) := X"10";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"10";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 106 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"10";
                        v_return(code*g_char_h + 2) := X"00";
                        v_return(code*g_char_h + 3) := X"10";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"10";
                        v_return(code*g_char_h + 6) := X"10";
                        v_return(code*g_char_h + 7) := X"70";
                    WHEN 107 =>
                        v_return(code*g_char_h + 0) := X"20";
                        v_return(code*g_char_h + 1) := X"20";
                        v_return(code*g_char_h + 2) := X"24";
                        v_return(code*g_char_h + 3) := X"38";
                        v_return(code*g_char_h + 4) := X"24";
                        v_return(code*g_char_h + 5) := X"24";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 108 =>
                        v_return(code*g_char_h + 0) := X"20";
                        v_return(code*g_char_h + 1) := X"20";
                        v_return(code*g_char_h + 2) := X"20";
                        v_return(code*g_char_h + 3) := X"20";
                        v_return(code*g_char_h + 4) := X"20";
                        v_return(code*g_char_h + 5) := X"38";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 109 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"63";
                        v_return(code*g_char_h + 3) := X"55";
                        v_return(code*g_char_h + 4) := X"49";
                        v_return(code*g_char_h + 5) := X"41";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 110 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"2E";
                        v_return(code*g_char_h + 3) := X"11";
                        v_return(code*g_char_h + 4) := X"11";
                        v_return(code*g_char_h + 5) := X"11";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 111 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"1C";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"1C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 112 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"3C";
                        v_return(code*g_char_h + 6) := X"20";
                        v_return(code*g_char_h + 7) := X"20";
                    WHEN 113 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"1E";
                        v_return(code*g_char_h + 3) := X"22";
                        v_return(code*g_char_h + 4) := X"22";
                        v_return(code*g_char_h + 5) := X"1E";
                        v_return(code*g_char_h + 6) := X"02";
                        v_return(code*g_char_h + 7) := X"02";
                    WHEN 114 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"2C";
                        v_return(code*g_char_h + 3) := X"12";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"10";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 115 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"3C";
                        v_return(code*g_char_h + 2) := X"22";
                        v_return(code*g_char_h + 3) := X"18";
                        v_return(code*g_char_h + 4) := X"44";
                        v_return(code*g_char_h + 5) := X"38";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 116 =>
                        v_return(code*g_char_h + 0) := X"10";
                        v_return(code*g_char_h + 1) := X"10";
                        v_return(code*g_char_h + 2) := X"38";
                        v_return(code*g_char_h + 3) := X"10";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"10";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 117 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"24";
                        v_return(code*g_char_h + 3) := X"24";
                        v_return(code*g_char_h + 4) := X"24";
                        v_return(code*g_char_h + 5) := X"18";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 118 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"14";
                        v_return(code*g_char_h + 3) := X"14";
                        v_return(code*g_char_h + 4) := X"14";
                        v_return(code*g_char_h + 5) := X"08";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 119 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"41";
                        v_return(code*g_char_h + 3) := X"49";
                        v_return(code*g_char_h + 4) := X"55";
                        v_return(code*g_char_h + 5) := X"63";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 120 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"24";
                        v_return(code*g_char_h + 3) := X"18";
                        v_return(code*g_char_h + 4) := X"18";
                        v_return(code*g_char_h + 5) := X"24";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 121 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"24";
                        v_return(code*g_char_h + 3) := X"24";
                        v_return(code*g_char_h + 4) := X"24";
                        v_return(code*g_char_h + 5) := X"3C";
                        v_return(code*g_char_h + 6) := X"04";
                        v_return(code*g_char_h + 7) := X"3C";
                    WHEN 122 =>
                        v_return(code*g_char_h + 0) := X"00";
                        v_return(code*g_char_h + 1) := X"00";
                        v_return(code*g_char_h + 2) := X"3C";
                        v_return(code*g_char_h + 3) := X"08";
                        v_return(code*g_char_h + 4) := X"10";
                        v_return(code*g_char_h + 5) := X"3C";
                        v_return(code*g_char_h + 6) := X"00";
                        v_return(code*g_char_h + 7) := X"00";
                    WHEN 123 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 124 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 125 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 126 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN 127 =>
                        v_return(code*g_char_h + 0) := "00000000";
                        v_return(code*g_char_h + 1) := "00000000";
                        v_return(code*g_char_h + 2) := "00000000";
                        v_return(code*g_char_h + 3) := "00000000";
                        v_return(code*g_char_h + 4) := "00000000";
                        v_return(code*g_char_h + 5) := "00000000";
                        v_return(code*g_char_h + 6) := "00000000";
                        v_return(code*g_char_h + 7) := "00000000";
                    WHEN OTHERS =>
                        NULL;
                END CASE;
            END LOOP;
        ELSE
            REPORT "character_ram: " &
                   integer'IMAGE(g_char_w) &
                   "x" &
                   integer'IMAGE(g_char_w) &
                   " characters, you're on your own - leaving character RAM empty, initialize it yourself"
                   SEVERITY warning;
        END IF;
        RETURN v_return;
    END FUNCTION;

    SIGNAL   r_char_arr : T_char_arr := f_init_char_arr;

BEGIN

    o_rd_data <= r_char_arr(to_integer(unsigned(i_rd_addr)));

    P_write : PROCESS(i_clk)
    BEGIN
        IF (rising_edge(i_clk)) THEN
            IF (i_wr_ena = '1') THEN
                r_char_arr(to_integer(unsigned(i_wr_addr))) <= i_wr_data;
            END IF;
        END IF;
    END PROCESS;

END ARCHITECTURE;
